ROM_RAWDATA_inst : ROM_RAWDATA PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		rden	 => rden_sig,
		q	 => q_sig
	);
